
module uart_rx_to_tx (

)



endmodule
